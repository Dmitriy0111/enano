`ifndef AHB_AGENT_PKG__SV
`define AHB_AGENT_PKG__SV

//  Package: ahb_agent_pkg
//
package ahb_agent_pkg;
    
    import uvm_pkg::*;

    `include "uvm_macros.svh"

    `include "ahb_item.sv"
    `include "ahb_agent_cfg.sv"
    
endpackage : ahb_agent_pkg

`endif // AHB_AGENT_PKG__SV
