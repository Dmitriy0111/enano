package uart_agent_pkg;

    import uvm_pkg::*;

    `include "uvm_macros.svh"
    `include "uart_item.sv"
    `include "uart_driver.sv"
    `include "uart_monitor.sv"
    `include "uart_agent_cfg.sv"
    `include "uart_item.sv"
    `include "uart_base_seq.sv"
    `include "uart_rand_seq.sv"
    `include "uart_sequencer.sv"
    `include "uart_subscriber.sv"
    `include "uart_agent.sv"

endpackage : uart_agent_pkg
