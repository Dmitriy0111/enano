module task_4;

    typedef struct{
        integer     ar[2];
    } ar_;

    ar_ pokr[$];

    initial
    begin
        $stop;
    end

endmodule : task_4
