package task_3_apb_pkg_ex;

    import      uvm_pkg::*;
    `include    "uvm_macros.svh"

    `include "task_3_apb_item_ex.sv"
    `include "task_3_apb_base_seq_ex.sv"
    `include "task_3_apb_rand_seq_ex.sv"
    `include "task_3_apb_sequencer_ex.sv"
    `include "task_3_apb_agent_cfg_ex.sv"
    `include "task_3_apb_master_ex.sv"
    `include "task_3_apb_monitor_ex.sv"
    `include "task_3_apb_agent_ex.sv"
    `include "task_3_apb_tb_env_ex.sv"
    `include "task_3_apb_base_test_ex.sv"
    `include "task_3_apb_run_item_test_ex.sv"

endpackage : task_3_apb_pkg_ex
