`ifndef APB_AGENT_PKG__SV
`define APB_AGENT_PKG__SV

//  Package: apb_agent_pkg
//
package apb_agent_pkg;
    
    import uvm_pkg::*;

    `include "uvm_macros.svh"

    `include "apb_item.sv"
    `include "apb_agent_cfg.sv"
    
endpackage : apb_agent_pkg

`endif // APB_AGENT_PKG__SV
