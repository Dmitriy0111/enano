//  Package: apb_test_pkg
//
package apb_test_pkg;
    // for UVM
    import uvm_pkg::*;
    
    import apb_agent_pkg::*;
    
    
    `include "uvm_macros.svh"
    `include "apb_env.sv"
    `include "apb_base_test.sv"
    `include "apb_run_item_test.sv"
    
endpackage : apb_test_pkg
