package uart_run_item_test_pkg;

    import uvm_pkg::*;

    import uart_agent_pkg::*;

    `include "uvm_macros.svh"
    `include "uart_env.sv"
    `include "uart_base_test.sv"
    `include "uart_run_item_test.sv"

endpackage : uart_run_item_test_pkg
