//  Package: axi_test_pkg
//
package axi_test_pkg;
    // for UVM
    import uvm_pkg::*;
    
    import axi_agent_pkg::*;
    
    `include "uvm_macros.svh"
    `include "axi_env.sv"
    `include "axi_base_test.sv"
    `include "axi_run_test.sv"
    
endpackage : axi_test_pkg
