//  Package: apb_agent_pkg
//
package apb_agent_pkg;
    // for UVM
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "apb_item.sv"
    `include "apb_base_seq.sv"
    `include "apb_rand_seq.sv"
    `include "apb_sequencer.sv"
    `include "apb_agent_cfg.sv"
    `include "apb_driver.sv"
    `include "apb_monitor.sv"
    `include "apb_agent.sv"
    
endpackage : apb_agent_pkg
